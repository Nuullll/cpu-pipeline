
module DataMemory(
    input clk,
    input rst_n,
    input [31:0] Address,
    input [31:0] Write_data,
    input MemRead,
    input MemWrite,

    output irqout,
    output reg [31:0] Read_data
);
    
    parameter RAM_SIZE = 512;
    parameter RAM_SIZE_BIT = 9;
    
    reg [31:0] RAM[RAM_SIZE - 1: 0];
    reg [31:0] TH,TL;
    reg [2:0]  TCON;
    reg        TCON_r1, TCON_r2;
    assign irqout = TCON[2];
    
    always @(*) 
    begin
        case(Address)
            32'h40000000: Read_data <= MemRead? TH: 32'd0;
            32'h40000004: Read_data <= MemRead? TL: 32'd0;
            32'h40000008: Read_data <= MemRead? {29'b0,TCON}: 32'd0;
            default: Read_data <= MemRead? RAM[Address[RAM_SIZE_BIT+1:2]]: 32'd0;
        endcase
    end
    
    always@(negedge rst_n or posedge clk) 
    begin
        if(~rst_n) begin
            TH <= 32'b0;
            TL <= 32'b0;
            TCON <= 3'b0;   
        end else begin
            TCON_r1 <= TCON[1];  
            TCON_r2 <= TCON_r1;
            if(TCON[0]) begin       //timer is enabled
                if(TL==32'hffffffff) begin
                    TL <= TH;
                    if(TCON[1]) TCON[2] <= 1'b1;        //irq is enabled
                end else TL <= TL + 1;
            end
            if(MemWrite) begin
                case(Address)
                    32'h40000000: TH <= Write_data;
                    32'h40000004: TL <= Write_data;
                    32'h40000008: TCON <= Write_data[2:0];      
                    default: ;
                endcase
            end
        end
    end
    

    always @(negedge rst_n or posedge clk)
        if (~rst_n) begin
            RAM[0] <= 32'h0000_0032; 
            RAM[1] <= 32'h0000_0043; 
            RAM[2] <= 32'h0000_00f6; 
            RAM[3] <= 32'h0000_00a8; 
            RAM[4] <= 32'h0000_0088; 
            RAM[5] <= 32'h0000_005a; 
            RAM[6] <= 32'h0000_0030; 
            RAM[7] <= 32'h0000_008d; 
            RAM[8] <= 32'h0000_0031; 
            RAM[9] <= 32'h0000_0031; 
            RAM[10] <= 32'h0000_0098; 
            RAM[11] <= 32'h0000_00a2; 
            RAM[12] <= 32'h0000_00e0; 
            RAM[13] <= 32'h0000_0037; 
            RAM[14] <= 32'h0000_0007; 
            RAM[15] <= 32'h0000_0034; 
            RAM[16] <= 32'h0000_002b; 
            RAM[17] <= 32'h0000_007e; 
            RAM[18] <= 32'h0000_0015; 
            RAM[19] <= 32'h0000_0016; 
            RAM[20] <= 32'h0000_0028; 
            RAM[21] <= 32'h0000_00ae; 
            RAM[22] <= 32'h0000_00d2; 
            RAM[23] <= 32'h0000_00a6; 
            RAM[24] <= 32'h0000_00ab; 
            RAM[25] <= 32'h0000_00f7; 
            RAM[26] <= 32'h0000_0015; 
            RAM[27] <= 32'h0000_0088; 
            RAM[28] <= 32'h0000_0009; 
            RAM[29] <= 32'h0000_00cf; 
            RAM[30] <= 32'h0000_004f; 
            RAM[31] <= 32'h0000_003c;
            RAM[32] <= 32'h0000_0000;
            RAM[33] <= 32'h0000_0000;
            RAM[34] <= 32'h0000_0000;
            RAM[35] <= 32'h0000_0000;
            RAM[36] <= 32'h0000_0000;
            RAM[37] <= 32'h0000_0000;
            RAM[38] <= 32'h0000_0000;
            RAM[39] <= 32'h0000_0000;
            RAM[40] <= 32'h0000_0000;
            RAM[41] <= 32'h0000_0000;
            RAM[42] <= 32'h0000_0000;
            RAM[43] <= 32'h0000_0000;
            RAM[44] <= 32'h0000_0000;
            RAM[45] <= 32'h0000_0000;
            RAM[46] <= 32'h0000_0000;
            RAM[47] <= 32'h0000_0000;
            RAM[48] <= 32'h0000_0000;
            RAM[49] <= 32'h0000_0000;
            RAM[50] <= 32'h0000_0000;
            RAM[51] <= 32'h0000_0000;
            RAM[52] <= 32'h0000_0000;
            RAM[53] <= 32'h0000_0000;
            RAM[54] <= 32'h0000_0000;
            RAM[55] <= 32'h0000_0000;
            RAM[56] <= 32'h0000_0000;
            RAM[57] <= 32'h0000_0000;
            RAM[58] <= 32'h0000_0000;
            RAM[59] <= 32'h0000_0000;
            RAM[60] <= 32'h0000_0000;
            RAM[61] <= 32'h0000_0000;
            RAM[62] <= 32'h0000_0000;
            RAM[63] <= 32'h0000_0000;
            RAM[64] <= 32'h0000_0000;
            RAM[65] <= 32'h0000_0000;
            RAM[66] <= 32'h0000_0000;
            RAM[67] <= 32'h0000_0000;
            RAM[68] <= 32'h0000_0000;
            RAM[69] <= 32'h0000_0000;
            RAM[70] <= 32'h0000_0000;
            RAM[71] <= 32'h0000_0000;
            RAM[72] <= 32'h0000_0000;
            RAM[73] <= 32'h0000_0000;
            RAM[74] <= 32'h0000_0000;
            RAM[75] <= 32'h0000_0000;
            RAM[76] <= 32'h0000_0000;
            RAM[77] <= 32'h0000_0000;
            RAM[78] <= 32'h0000_0000;
            RAM[79] <= 32'h0000_0000;
            RAM[80] <= 32'h0000_0000;
            RAM[81] <= 32'h0000_0000;
            RAM[82] <= 32'h0000_0000;
            RAM[83] <= 32'h0000_0000;
            RAM[84] <= 32'h0000_0000;
            RAM[85] <= 32'h0000_0000;
            RAM[86] <= 32'h0000_0000;
            RAM[87] <= 32'h0000_0000;
            RAM[88] <= 32'h0000_0000;
            RAM[89] <= 32'h0000_0000;
            RAM[90] <= 32'h0000_0000;
            RAM[91] <= 32'h0000_0000;
            RAM[92] <= 32'h0000_0000;
            RAM[93] <= 32'h0000_0000;
            RAM[94] <= 32'h0000_0000;
            RAM[95] <= 32'h0000_0000;
            RAM[96] <= 32'h0000_0000;
            RAM[97] <= 32'h0000_0000;
            RAM[98] <= 32'h0000_0000;
            RAM[99] <= 32'h0000_0000;
            RAM[100] <= 32'h0000_0000;
            RAM[101] <= 32'h0000_0000;
            RAM[102] <= 32'h0000_0000;
            RAM[103] <= 32'h0000_0000;
            RAM[104] <= 32'h0000_0000;
            RAM[105] <= 32'h0000_0000;
            RAM[106] <= 32'h0000_0000;
            RAM[107] <= 32'h0000_0000;
            RAM[108] <= 32'h0000_0000;
            RAM[109] <= 32'h0000_0000;
            RAM[110] <= 32'h0000_0000;
            RAM[111] <= 32'h0000_0000;
            RAM[112] <= 32'h0000_0000;
            RAM[113] <= 32'h0000_0000;
            RAM[114] <= 32'h0000_0000;
            RAM[115] <= 32'h0000_0000;
            RAM[116] <= 32'h0000_0000;
            RAM[117] <= 32'h0000_0000;
            RAM[118] <= 32'h0000_0000;
            RAM[119] <= 32'h0000_0000;
            RAM[120] <= 32'h0000_0000;
            RAM[121] <= 32'h0000_0000;
            RAM[122] <= 32'h0000_0000;
            RAM[123] <= 32'h0000_0000;
            RAM[124] <= 32'h0000_0000;
            RAM[125] <= 32'h0000_0000;
            RAM[126] <= 32'h0000_0000;
            RAM[127] <= 32'h0000_0000;
            RAM[128] <= 32'h0000_0000;
            RAM[129] <= 32'h0000_0000;
            RAM[130] <= 32'h0000_0000;
            RAM[131] <= 32'h0000_0000;
            RAM[132] <= 32'h0000_0000;
            RAM[133] <= 32'h0000_0000;
            RAM[134] <= 32'h0000_0000;
            RAM[135] <= 32'h0000_0000;
            RAM[136] <= 32'h0000_0000;
            RAM[137] <= 32'h0000_0000;
            RAM[138] <= 32'h0000_0000;
            RAM[139] <= 32'h0000_0000;
            RAM[140] <= 32'h0000_0000;
            RAM[141] <= 32'h0000_0000;
            RAM[142] <= 32'h0000_0000;
            RAM[143] <= 32'h0000_0000;
            RAM[144] <= 32'h0000_0000;
            RAM[145] <= 32'h0000_0000;
            RAM[146] <= 32'h0000_0000;
            RAM[147] <= 32'h0000_0000;
            RAM[148] <= 32'h0000_0000;
            RAM[149] <= 32'h0000_0000;
            RAM[150] <= 32'h0000_0000;
            RAM[151] <= 32'h0000_0000;
            RAM[152] <= 32'h0000_0000;
            RAM[153] <= 32'h0000_0000;
            RAM[154] <= 32'h0000_0000;
            RAM[155] <= 32'h0000_0000;
            RAM[156] <= 32'h0000_0000;
            RAM[157] <= 32'h0000_0000;
            RAM[158] <= 32'h0000_0000;
            RAM[159] <= 32'h0000_0000;
            RAM[160] <= 32'h0000_0000;
            RAM[161] <= 32'h0000_0000;
            RAM[162] <= 32'h0000_0000;
            RAM[163] <= 32'h0000_0000;
            RAM[164] <= 32'h0000_0000;
            RAM[165] <= 32'h0000_0000;
            RAM[166] <= 32'h0000_0000;
            RAM[167] <= 32'h0000_0000;
            RAM[168] <= 32'h0000_0000;
            RAM[169] <= 32'h0000_0000;
            RAM[170] <= 32'h0000_0000;
            RAM[171] <= 32'h0000_0000;
            RAM[172] <= 32'h0000_0000;
            RAM[173] <= 32'h0000_0000;
            RAM[174] <= 32'h0000_0000;
            RAM[175] <= 32'h0000_0000;
            RAM[176] <= 32'h0000_0000;
            RAM[177] <= 32'h0000_0000;
            RAM[178] <= 32'h0000_0000;
            RAM[179] <= 32'h0000_0000;
            RAM[180] <= 32'h0000_0000;
            RAM[181] <= 32'h0000_0000;
            RAM[182] <= 32'h0000_0000;
            RAM[183] <= 32'h0000_0000;
            RAM[184] <= 32'h0000_0000;
            RAM[185] <= 32'h0000_0000;
            RAM[186] <= 32'h0000_0000;
            RAM[187] <= 32'h0000_0000;
            RAM[188] <= 32'h0000_0000;
            RAM[189] <= 32'h0000_0000;
            RAM[190] <= 32'h0000_0000;
            RAM[191] <= 32'h0000_0000;
            RAM[192] <= 32'h0000_0000;
            RAM[193] <= 32'h0000_0000;
            RAM[194] <= 32'h0000_0000;
            RAM[195] <= 32'h0000_0000;
            RAM[196] <= 32'h0000_0000;
            RAM[197] <= 32'h0000_0000;
            RAM[198] <= 32'h0000_0000;
            RAM[199] <= 32'h0000_0000;
            RAM[200] <= 32'h0000_0000;
            RAM[201] <= 32'h0000_0000;
            RAM[202] <= 32'h0000_0000;
            RAM[203] <= 32'h0000_0000;
            RAM[204] <= 32'h0000_0000;
            RAM[205] <= 32'h0000_0000;
            RAM[206] <= 32'h0000_0000;
            RAM[207] <= 32'h0000_0000;
            RAM[208] <= 32'h0000_0000;
            RAM[209] <= 32'h0000_0000;
            RAM[210] <= 32'h0000_0000;
            RAM[211] <= 32'h0000_0000;
            RAM[212] <= 32'h0000_0000;
            RAM[213] <= 32'h0000_0000;
            RAM[214] <= 32'h0000_0000;
            RAM[215] <= 32'h0000_0000;
            RAM[216] <= 32'h0000_0000;
            RAM[217] <= 32'h0000_0000;
            RAM[218] <= 32'h0000_0000;
            RAM[219] <= 32'h0000_0000;
            RAM[220] <= 32'h0000_0000;
            RAM[221] <= 32'h0000_0000;
            RAM[222] <= 32'h0000_0000;
            RAM[223] <= 32'h0000_0000;
            RAM[224] <= 32'h0000_0000;
            RAM[225] <= 32'h0000_0000;
            RAM[226] <= 32'h0000_0000;
            RAM[227] <= 32'h0000_0000;
            RAM[228] <= 32'h0000_0000;
            RAM[229] <= 32'h0000_0000;
            RAM[230] <= 32'h0000_0000;
            RAM[231] <= 32'h0000_0000;
            RAM[232] <= 32'h0000_0000;
            RAM[233] <= 32'h0000_0000;
            RAM[234] <= 32'h0000_0000;
            RAM[235] <= 32'h0000_0000;
            RAM[236] <= 32'h0000_0000;
            RAM[237] <= 32'h0000_0000;
            RAM[238] <= 32'h0000_0000;
            RAM[239] <= 32'h0000_0000;
            RAM[240] <= 32'h0000_0000;
            RAM[241] <= 32'h0000_0000;
            RAM[242] <= 32'h0000_0000;
            RAM[243] <= 32'h0000_0000;
            RAM[244] <= 32'h0000_0000;
            RAM[245] <= 32'h0000_0000;
            RAM[246] <= 32'h0000_0000;
            RAM[247] <= 32'h0000_0000;
            RAM[248] <= 32'h0000_0000;
            RAM[249] <= 32'h0000_0000;
            RAM[250] <= 32'h0000_0000;
            RAM[251] <= 32'h0000_0000;
            RAM[252] <= 32'h0000_0000;
            RAM[253] <= 32'h0000_0000;
            RAM[254] <= 32'h0000_0000;
            RAM[255] <= 32'h0000_0000;
            RAM[256] <= 32'h0000_0063; 
            RAM[257] <= 32'h0000_007c; 
            RAM[258] <= 32'h0000_0077; 
            RAM[259] <= 32'h0000_007b; 
            RAM[260] <= 32'h0000_00f2; 
            RAM[261] <= 32'h0000_006b; 
            RAM[262] <= 32'h0000_006f; 
            RAM[263] <= 32'h0000_00c5; 
            RAM[264] <= 32'h0000_0030; 
            RAM[265] <= 32'h0000_0001; 
            RAM[266] <= 32'h0000_0067; 
            RAM[267] <= 32'h0000_002b; 
            RAM[268] <= 32'h0000_00fe; 
            RAM[269] <= 32'h0000_00d7; 
            RAM[270] <= 32'h0000_00ab; 
            RAM[271] <= 32'h0000_0076; 
            RAM[272] <= 32'h0000_00ca; 
            RAM[273] <= 32'h0000_0082; 
            RAM[274] <= 32'h0000_00c9; 
            RAM[275] <= 32'h0000_007d; 
            RAM[276] <= 32'h0000_00fa; 
            RAM[277] <= 32'h0000_0059; 
            RAM[278] <= 32'h0000_0047; 
            RAM[279] <= 32'h0000_00f0; 
            RAM[280] <= 32'h0000_00ad; 
            RAM[281] <= 32'h0000_00d4; 
            RAM[282] <= 32'h0000_00a2; 
            RAM[283] <= 32'h0000_00af; 
            RAM[284] <= 32'h0000_009c; 
            RAM[285] <= 32'h0000_00a4; 
            RAM[286] <= 32'h0000_0072; 
            RAM[287] <= 32'h0000_00c0; 
            RAM[288] <= 32'h0000_00b7; 
            RAM[289] <= 32'h0000_00fd; 
            RAM[290] <= 32'h0000_0093; 
            RAM[291] <= 32'h0000_0026; 
            RAM[292] <= 32'h0000_0036; 
            RAM[293] <= 32'h0000_003f; 
            RAM[294] <= 32'h0000_00f7; 
            RAM[295] <= 32'h0000_00cc; 
            RAM[296] <= 32'h0000_0034; 
            RAM[297] <= 32'h0000_00a5; 
            RAM[298] <= 32'h0000_00e5; 
            RAM[299] <= 32'h0000_00f1; 
            RAM[300] <= 32'h0000_0071; 
            RAM[301] <= 32'h0000_00d8; 
            RAM[302] <= 32'h0000_0031; 
            RAM[303] <= 32'h0000_0015; 
            RAM[304] <= 32'h0000_0004; 
            RAM[305] <= 32'h0000_00c7; 
            RAM[306] <= 32'h0000_0023; 
            RAM[307] <= 32'h0000_00c3; 
            RAM[308] <= 32'h0000_0018; 
            RAM[309] <= 32'h0000_0096; 
            RAM[310] <= 32'h0000_0005; 
            RAM[311] <= 32'h0000_009a; 
            RAM[312] <= 32'h0000_0007; 
            RAM[313] <= 32'h0000_0012; 
            RAM[314] <= 32'h0000_0080; 
            RAM[315] <= 32'h0000_00e2; 
            RAM[316] <= 32'h0000_00eb; 
            RAM[317] <= 32'h0000_0027; 
            RAM[318] <= 32'h0000_00b2; 
            RAM[319] <= 32'h0000_0075; 
            RAM[320] <= 32'h0000_0009; 
            RAM[321] <= 32'h0000_0083; 
            RAM[322] <= 32'h0000_002c; 
            RAM[323] <= 32'h0000_001a; 
            RAM[324] <= 32'h0000_001b; 
            RAM[325] <= 32'h0000_006e; 
            RAM[326] <= 32'h0000_005a; 
            RAM[327] <= 32'h0000_00a0; 
            RAM[328] <= 32'h0000_0052; 
            RAM[329] <= 32'h0000_003b; 
            RAM[330] <= 32'h0000_00d6; 
            RAM[331] <= 32'h0000_00b3; 
            RAM[332] <= 32'h0000_0029; 
            RAM[333] <= 32'h0000_00e3; 
            RAM[334] <= 32'h0000_002f; 
            RAM[335] <= 32'h0000_0084; 
            RAM[336] <= 32'h0000_0053; 
            RAM[337] <= 32'h0000_00d1; 
            RAM[338] <= 32'h0000_0000; 
            RAM[339] <= 32'h0000_00ed; 
            RAM[340] <= 32'h0000_0020; 
            RAM[341] <= 32'h0000_00fc; 
            RAM[342] <= 32'h0000_00b1; 
            RAM[343] <= 32'h0000_005b; 
            RAM[344] <= 32'h0000_006a; 
            RAM[345] <= 32'h0000_00cb; 
            RAM[346] <= 32'h0000_00be; 
            RAM[347] <= 32'h0000_0039; 
            RAM[348] <= 32'h0000_004a; 
            RAM[349] <= 32'h0000_004c; 
            RAM[350] <= 32'h0000_0058; 
            RAM[351] <= 32'h0000_00cf; 
            RAM[352] <= 32'h0000_00d0; 
            RAM[353] <= 32'h0000_00ef; 
            RAM[354] <= 32'h0000_00aa; 
            RAM[355] <= 32'h0000_00fb; 
            RAM[356] <= 32'h0000_0043; 
            RAM[357] <= 32'h0000_004d; 
            RAM[358] <= 32'h0000_0033; 
            RAM[359] <= 32'h0000_0085; 
            RAM[360] <= 32'h0000_0045; 
            RAM[361] <= 32'h0000_00f9; 
            RAM[362] <= 32'h0000_0002; 
            RAM[363] <= 32'h0000_007f; 
            RAM[364] <= 32'h0000_0050; 
            RAM[365] <= 32'h0000_003c; 
            RAM[366] <= 32'h0000_009f; 
            RAM[367] <= 32'h0000_00a8; 
            RAM[368] <= 32'h0000_0051; 
            RAM[369] <= 32'h0000_00a3; 
            RAM[370] <= 32'h0000_0040; 
            RAM[371] <= 32'h0000_008f; 
            RAM[372] <= 32'h0000_0092; 
            RAM[373] <= 32'h0000_009d; 
            RAM[374] <= 32'h0000_0038; 
            RAM[375] <= 32'h0000_00f5; 
            RAM[376] <= 32'h0000_00bc; 
            RAM[377] <= 32'h0000_00b6; 
            RAM[378] <= 32'h0000_00da; 
            RAM[379] <= 32'h0000_0021; 
            RAM[380] <= 32'h0000_0010; 
            RAM[381] <= 32'h0000_00ff; 
            RAM[382] <= 32'h0000_00f3; 
            RAM[383] <= 32'h0000_00d2; 
            RAM[384] <= 32'h0000_00cd; 
            RAM[385] <= 32'h0000_000c; 
            RAM[386] <= 32'h0000_0013; 
            RAM[387] <= 32'h0000_00ec; 
            RAM[388] <= 32'h0000_005f; 
            RAM[389] <= 32'h0000_0097; 
            RAM[390] <= 32'h0000_0044; 
            RAM[391] <= 32'h0000_0017; 
            RAM[392] <= 32'h0000_00c4; 
            RAM[393] <= 32'h0000_00a7; 
            RAM[394] <= 32'h0000_007e; 
            RAM[395] <= 32'h0000_003d; 
            RAM[396] <= 32'h0000_0064; 
            RAM[397] <= 32'h0000_005d; 
            RAM[398] <= 32'h0000_0019; 
            RAM[399] <= 32'h0000_0073; 
            RAM[400] <= 32'h0000_0060; 
            RAM[401] <= 32'h0000_0081; 
            RAM[402] <= 32'h0000_004f; 
            RAM[403] <= 32'h0000_00dc; 
            RAM[404] <= 32'h0000_0022; 
            RAM[405] <= 32'h0000_002a; 
            RAM[406] <= 32'h0000_0090; 
            RAM[407] <= 32'h0000_0088; 
            RAM[408] <= 32'h0000_0046; 
            RAM[409] <= 32'h0000_00ee; 
            RAM[410] <= 32'h0000_00b8; 
            RAM[411] <= 32'h0000_0014; 
            RAM[412] <= 32'h0000_00de; 
            RAM[413] <= 32'h0000_005e; 
            RAM[414] <= 32'h0000_000b; 
            RAM[415] <= 32'h0000_00db; 
            RAM[416] <= 32'h0000_00e0; 
            RAM[417] <= 32'h0000_0032; 
            RAM[418] <= 32'h0000_003a; 
            RAM[419] <= 32'h0000_000a; 
            RAM[420] <= 32'h0000_0049; 
            RAM[421] <= 32'h0000_0006; 
            RAM[422] <= 32'h0000_0024; 
            RAM[423] <= 32'h0000_005c; 
            RAM[424] <= 32'h0000_00c2; 
            RAM[425] <= 32'h0000_00d3; 
            RAM[426] <= 32'h0000_00ac; 
            RAM[427] <= 32'h0000_0062; 
            RAM[428] <= 32'h0000_0091; 
            RAM[429] <= 32'h0000_0095; 
            RAM[430] <= 32'h0000_00e4; 
            RAM[431] <= 32'h0000_0079; 
            RAM[432] <= 32'h0000_00e7; 
            RAM[433] <= 32'h0000_00c8; 
            RAM[434] <= 32'h0000_0037; 
            RAM[435] <= 32'h0000_006d; 
            RAM[436] <= 32'h0000_008d; 
            RAM[437] <= 32'h0000_00d5; 
            RAM[438] <= 32'h0000_004e; 
            RAM[439] <= 32'h0000_00a9; 
            RAM[440] <= 32'h0000_006c; 
            RAM[441] <= 32'h0000_0056; 
            RAM[442] <= 32'h0000_00f4; 
            RAM[443] <= 32'h0000_00ea; 
            RAM[444] <= 32'h0000_0065; 
            RAM[445] <= 32'h0000_007a; 
            RAM[446] <= 32'h0000_00ae; 
            RAM[447] <= 32'h0000_0008; 
            RAM[448] <= 32'h0000_00ba; 
            RAM[449] <= 32'h0000_0078; 
            RAM[450] <= 32'h0000_0025; 
            RAM[451] <= 32'h0000_002e; 
            RAM[452] <= 32'h0000_001c; 
            RAM[453] <= 32'h0000_00a6; 
            RAM[454] <= 32'h0000_00b4; 
            RAM[455] <= 32'h0000_00c6; 
            RAM[456] <= 32'h0000_00e8; 
            RAM[457] <= 32'h0000_00dd; 
            RAM[458] <= 32'h0000_0074; 
            RAM[459] <= 32'h0000_001f; 
            RAM[460] <= 32'h0000_004b; 
            RAM[461] <= 32'h0000_00bd; 
            RAM[462] <= 32'h0000_008b; 
            RAM[463] <= 32'h0000_008a; 
            RAM[464] <= 32'h0000_0070; 
            RAM[465] <= 32'h0000_003e; 
            RAM[466] <= 32'h0000_00b5; 
            RAM[467] <= 32'h0000_0066; 
            RAM[468] <= 32'h0000_0048; 
            RAM[469] <= 32'h0000_0003; 
            RAM[470] <= 32'h0000_00f6; 
            RAM[471] <= 32'h0000_000e; 
            RAM[472] <= 32'h0000_0061; 
            RAM[473] <= 32'h0000_0035; 
            RAM[474] <= 32'h0000_0057; 
            RAM[475] <= 32'h0000_00b9; 
            RAM[476] <= 32'h0000_0086; 
            RAM[477] <= 32'h0000_00c1; 
            RAM[478] <= 32'h0000_001d; 
            RAM[479] <= 32'h0000_009e; 
            RAM[480] <= 32'h0000_00e1; 
            RAM[481] <= 32'h0000_00f8; 
            RAM[482] <= 32'h0000_0098; 
            RAM[483] <= 32'h0000_0011; 
            RAM[484] <= 32'h0000_0069; 
            RAM[485] <= 32'h0000_00d9; 
            RAM[486] <= 32'h0000_008e; 
            RAM[487] <= 32'h0000_0094; 
            RAM[488] <= 32'h0000_009b; 
            RAM[489] <= 32'h0000_001e; 
            RAM[490] <= 32'h0000_0087; 
            RAM[491] <= 32'h0000_00e9; 
            RAM[492] <= 32'h0000_00ce; 
            RAM[493] <= 32'h0000_0055; 
            RAM[494] <= 32'h0000_0028; 
            RAM[495] <= 32'h0000_00df; 
            RAM[496] <= 32'h0000_008c; 
            RAM[497] <= 32'h0000_00a1; 
            RAM[498] <= 32'h0000_0089; 
            RAM[499] <= 32'h0000_000d; 
            RAM[500] <= 32'h0000_00bf; 
            RAM[501] <= 32'h0000_00e6; 
            RAM[502] <= 32'h0000_0042; 
            RAM[503] <= 32'h0000_0068; 
            RAM[504] <= 32'h0000_0041; 
            RAM[505] <= 32'h0000_0099; 
            RAM[506] <= 32'h0000_002d; 
            RAM[507] <= 32'h0000_000f; 
            RAM[508] <= 32'h0000_00b0; 
            RAM[509] <= 32'h0000_0054; 
            RAM[510] <= 32'h0000_00bb; 
            RAM[511] <= 32'h0000_0016;
        end else if (MemWrite && Address[RAM_SIZE_BIT+1:2] < RAM_SIZE) begin 
            RAM[Address[RAM_SIZE_BIT+1:2]] <= Write_data;
        end     

            
endmodule
